//write a module which acts like an inverter.
module top_module( input in, output out );
	assign out = ~in;
endmodule
