//write a code for simple wire declaration such that the input is 
//driven as the output one
module test_01(input in , output out);
	assign out = in ; //already in verilog the output variable is wire type
endmodule 
