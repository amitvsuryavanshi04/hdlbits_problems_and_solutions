//create a module that implements and gate 
module top_module( 
    input a, 
    input b, 
    output out );
	assign out = a & b;
endmodule
