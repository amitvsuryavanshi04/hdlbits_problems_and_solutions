// code which passes only value zero..... 

module top_module(
    output zero
);// Module body starts after semicolon
    assign zero = 1'b0;
	
endmodule

//write a code which passes value as only one 
module top_module_one(output one);
	assign one = 1'b1;
endmodule 

