/*
Quesiton:
implement a circuit which does following thing 
in <------------------------> out
*/

module top_module (
    input in,
    output out);
assign out = in ;
endmodule
