/*
Question:
You are provided with a BCD one-digit adder named bcd_fadd that 
adds two BCD digits and carry-in, and produces a sum and carry-out.

module bcd_fadd (
    input [3:0] a,
    input [3:0] b,
    input     cin,
    output   cout,
    output [3:0] sum );

Instantiate 100 copies of bcd_fadd to create a 100-digit BCD
 ripple-carry adder. Your adder should add two 100-digit BCD
  numbers (packed into 400-bit vectors) and a carry-in to 
  produce a 100-digit sum and carry out. 
*/
//solution
module top_module( 
    input [399:0] a, b,
    input cin,
    output cout,
    output [399:0] sum );
    wire[99:0] cout_wires;
    genvar gv;
    
    generate
        bcd_fadd(a[3:0], b[3:0], cin, cout_wires[0],sum[3:0]);
        for (gv=4; gv<400; gv=gv+4) begin: bcd_adder_instances
            bcd_fadd bcd_adder(a[gv+3:gv], b[gv+3:gv], cout_wires[gv/4-1],cout_wires[gv/4],sum[gv+3:gv]);
        end
    endgenerate
    
    assign cout = cout_wires[99];

endmodule
