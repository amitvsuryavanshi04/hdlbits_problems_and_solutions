/*
Quesiton:
implement the below circuit:
    ----------out
    |
    |
    |
  -----
   ---
    -

*/

//solution
module top_module(output out);
    assign out = 1'b0; //assign 1'b0 for the GND
endmodule
